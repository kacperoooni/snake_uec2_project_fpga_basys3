`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.09.2020 19:06:09
// Design Name: 
// Module Name: menu_display
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module key_debouncer(
	input wire clk,
	input wire [15:0] vcount, hcount,
	output wire vsync_in,hsync_in,hsync_out,vsync_out,
	input wire rx_empty,
	input wire [7:0] r_data,
	output reg [7:0] r_data_debug,
	output reg [7:0] key_data 
    );
    
  localparam
  INIT = 0,
  KEY_PRESSED = 1,
  KEY_RELASED = 2;
  
  reg [3:0] state, state_nxt;
  reg [7:0] key_data_nxt;
//  assign r_data_debug = key_data;  
    
 always@*
 	begin
    if(rx_empty == 0)
    	begin 
    		key_data_nxt = r_data;
    		r_data_debug = 8'hFF;
    	end	
    else 
    	begin
    		key_data_nxt = 8'b0;
    	end	
	end
   
 always@(posedge clk)
  begin
  	key_data = key_data_nxt;
  end	
    
    
    
endmodule
