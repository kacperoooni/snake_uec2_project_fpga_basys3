//Listing 8.4




//MODUL ZAIMPORTOWANY Z CWICZENIA NR 6 - UEC2
module uart
   #( // Default setting:
      // 9.600 baud, 8 data bits, 1 stop bit, 2^2 FIFO
      parameter DBIT = 8,     // # data bits
                SB_TICK = 16, // # ticks for stop bits, 16/24/32
                              // for 1/1.5/2 stop bits
                DVSR = 65000000/(16*9600),//DVSR = 326,   // baud rate divisor
                              // DVSR = 50M/(16*baud rate)
                DVSR_BIT = 9, // # bits of DVSR
                FIFO_W = 1    // # addr bits of FIFO
                              // # words in FIFO=2^FIFO_W
   )
   (
    input wire clk, reset,
    input wire  rx, //rd_uart, wr_uart,
  //  input wire [7:0] w_data,
    output wire  tx, rx_empty,
    output wire [7:0] r_data,
    output reg [7:0] word,
    output wire [7:0] led
   );

  
   // signal declaration
   wire tick, rx_done_tick, tx_done_tick;
   wire tx_empty, tx_fifo_not_empty;
   wire [7:0] tx_fifo_out, rx_data_out;
   wire [7:0] w_data;
   reg rd_uart, rd_uart_nxt;
  // wire [7:0] r_data;
   reg [7:0] word_nxt;
   assign w_data = 0;

   //body
   mod_m_counter #(.M(DVSR), .N(DVSR_BIT)) baud_gen_unit
      (.clk(clk), .reset(reset), .q(), .max_tick(tick));

   uart_rx #(.DBIT(DBIT), .SB_TICK(SB_TICK)) uart_rx_unit
      (.clk(clk), .reset(reset), .rx(rx), .s_tick(tick),
       .rx_done_tick(rx_done_tick), .dout(rx_data_out));

   fifo #(.B(DBIT), .W(FIFO_W)) fifo_rx_unit
      (.clk(clk), .reset(reset), .rd(rd_uart),
       .wr(rx_done_tick), .w_data(rx_data_out),
       .empty(rx_empty), .full(), .r_data(r_data));

   fifo #(.B(DBIT), .W(FIFO_W)) fifo_tx_unit
      (.clk(clk), .reset(reset), .rd(tx_done_tick),
       .wr(wr_uart), .w_data(w_data), .empty(tx_empty),
       .full(tx_full), .r_data(tx_fifo_out));

   uart_tx #(.DBIT(DBIT), .SB_TICK(SB_TICK)) uart_tx_unit
      (.clk(clk), .reset(reset), .tx_start(tx_fifo_not_empty),
       .s_tick(tick), .din(tx_fifo_out),
       .tx_done_tick(tx_done_tick), .tx(tx));

   assign tx_fifo_not_empty = ~tx_empty;
   
    always@(*)
    begin
    if((~rx_empty) && (rd_uart == 0))
        begin
        word_nxt = r_data;
        rd_uart_nxt = 1;
        end
    else if(reset)
    		begin
    		word_nxt = 0;
    		rd_uart_nxt = 0;
    		end   
    else
        begin
        word_nxt = word;
        rd_uart_nxt = 0;
        end    
    end
    
    always@(posedge clk)
    begin
    rd_uart <= rd_uart_nxt;
    word <= word_nxt;
    end
    assign led = word;
    

endmodule