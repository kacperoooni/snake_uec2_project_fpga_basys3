`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12.08.2020 23:42:23
// Design Name: 
// Module Name: rect_controller
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module rect_controller(
    output reg [31:0] rect_read_out,
    output reg [35:0] rect_write,
    output reg [15:0] score_out,
    output reg game_over,
    input wire [3:0] rect_read_in,
    input wire clk,
		input wire [7:0] key,
		input wire rst,
		input wire [7:0] r_data,
		input wire menu_interrupt, game_start,
		input wire [1:0] difficulty_level_in,
		input wire game_restart
		
		
	
	//DEBUG
	//	output reg [3:0] an,  // enable 1-out-of-4 asserted low
  //  output reg [6:0] sseg, // led segments
	//	input wire [4:0] debug_keys,
	//	input wire [15:0] iterator_debug 
	
	
    );
    wire [2:0] difficulty_level;
    assign difficulty_level = difficulty_level_in + 1;
   localparam 
      GRID_SIZE_X = 32,
      GRID_SIZE_Y = 24,
      RECT_SIZE_X = (1024/GRID_SIZE_X),
      RECT_SIZE_Y = (768/GRID_SIZE_Y),
      NULL = 4'b0000,
      SNAKE = 4'b0001,
      ROCK = 4'b0010,
      SNACK = 4'b0100;
   
   localparam
   	WAIT_FOR_START = 5'd0, //states
		INIT = 5'd1,
		SNAKE_MOVING = 5'd2,
		SNAKE_GROW = 5'd3,
		RESET = 5'd4,
		GAME_OVER = 5'd5,
		SNAKE_DRAWING = 5'd6,
		COLLISION_READ = 5'd7,
		COLLISION_CHECK = 5'd8,
		SNACK_GENERATE = 5'd9,
		SNACK_CHECK_READ = 5'd10,
		SNACK_CHECK_WRITE = 5'd11,
		MENU_INTERRUPT = 5'd12;
   
   localparam //keys
    UP = 8'h38,
    DOWN = 8'h32,
    LEFT = 8'h34,
    RIGHT = 8'h36,
    UP_RIGHT = 8'h39,
    UP_LEFT = 8'h37,
    DOWN_RIGHT = 8'h33,
    DOWN_LEFT = 8'h31,
    MIDDLE = 8'h35;
	
	
	localparam 
	SNAKE_REG_SIZE = 127,//+1
	//DIFFICULTY = 3,
	SNAKE_TURBO = 10000000; 
	
   
   reg [31:0] rect_read_out_nxt;
   reg [15:0] rect_read_x_nxt, rect_read_y_nxt;
   reg [4:0]  state;
   reg [4:0]  state_nxt;
   reg [35:0] rect_write_nxt;
   reg [31:0] snake_register [SNAKE_REG_SIZE:0];
   reg [31:0] snake_register_nxt [SNAKE_REG_SIZE:0];
   
   reg [15:0] score_nxt;
   reg [31:0] i; //intertor for smth
   reg [15:0] snake_writer_iterator, snake_writer_iterator_nxt; //interator for writing snake rects
   reg [31:0] snake_moving_iterator,snake_moving_iterator_nxt; //interator for moving period of snake
   
   

   reg [15:0] snake_size, snake_size_nxt;
   reg [31:0] previous_read_rect;
   reg [4:0] snack_gen_reg_y, snack_gen_reg_y_nxt, snack_gen_reg_x, snack_gen_reg_x_nxt;
   reg [31:0] snake_speed, snake_speed_nxt;
   reg game_over_nxt;
   
   
   
   
   
  //{rect_write_x,rect_write_y,rect_write_function} = rect_write;
   always@(*)
     begin
				state_nxt = WAIT_FOR_START;
				snake_moving_iterator_nxt = snake_moving_iterator + 1;
				snake_writer_iterator_nxt = snake_writer_iterator;
				snake_size_nxt = snake_size;
				rect_write_nxt = rect_write; //WARNING!! CAN CAUSE UNEXPECTED WRITE TO MEMORY
				snack_gen_reg_y_nxt = snack_gen_reg_y;
				snack_gen_reg_x_nxt = snack_gen_reg_x;
				rect_read_out_nxt = rect_read_out;
				snake_speed_nxt = snake_speed;
				score_nxt = score_out;
				game_over_nxt = game_over;
				for(i = 0; i <= SNAKE_REG_SIZE; i=i+1)
					begin
						snake_register_nxt[i] = snake_register[i];
					end


				case(state)
					WAIT_FOR_START:
						begin
							if(game_start == 1) state_nxt = INIT;
							else state_nxt = WAIT_FOR_START;
							game_over_nxt = 0; 
						end	
					INIT:
						begin
							for(i = 0; i <= SNAKE_REG_SIZE; i=i+1)
							begin
								snake_register_nxt[i] = 0;
							end
							snake_register_nxt[0] = {16'd15,16'd15};
							snake_register_nxt[1] = {16'd16,16'd15};
							snake_register_nxt[2] = {16'd17,16'd15};
							snake_register_nxt[3] = {16'd18,16'd15};
							snake_size_nxt = 3; // with 0
							snake_writer_iterator_nxt = 0;
							snake_moving_iterator_nxt = 0;
							snake_speed_nxt = 50000000;
							state_nxt = SNAKE_MOVING;
							score_nxt = 0;
							game_over_nxt = 0;
						end

					SNAKE_MOVING:
						begin
							state_nxt = COLLISION_READ;
							snake_moving_iterator_nxt = 0;
							for(i = 0; i < SNAKE_REG_SIZE; i=i+1)
							begin
								snake_register_nxt[i+1] = snake_register[i]; //shift snake stack
							end
							case(key)
								DOWN:
								begin
									snake_register_nxt[0] = {snake_register[0][31:16],snake_register[0][15:0]+16'd1};
								end
								LEFT:
								begin
									snake_register_nxt[0] = {snake_register[0][31:16]-16'd1,snake_register[0][15:0]};
								end
								RIGHT:
								begin
									snake_register_nxt[0] = {snake_register[0][31:16]+16'd1,snake_register[0][15:0]};
								end
								UP:
								begin
									snake_register_nxt[0] = {snake_register[0][31:16],snake_register[0][15:0]-16'd1};
								end
								DOWN_RIGHT:
								begin
									snake_register_nxt[0] = {snake_register[0][31:16]+16'd1,snake_register[0][15:0]+16'd1};
								end
								DOWN_LEFT:
								begin
									snake_register_nxt[0] = {snake_register[0][31:16]-16'd1,snake_register[0][15:0]+16'd1};
								end
								UP_RIGHT:
								begin
									snake_register_nxt[0] = {snake_register[0][31:16]+16'd1,snake_register[0][15:0]-16'd1};
								end
								UP_LEFT:
								begin
									snake_register_nxt[0] = {snake_register[0][31:16]-16'd1,snake_register[0][15:0]-16'd1};
								end
								default: begin end
							endcase
						end

					SNAKE_DRAWING:
						begin
							if(snake_moving_iterator == snake_speed)	state_nxt = SNAKE_MOVING;
							else if(menu_interrupt == 1) state_nxt = MENU_INTERRUPT;
							else state_nxt = SNAKE_DRAWING;

							if(snake_register[snake_writer_iterator] != 0)
							rect_write_nxt = {snake_register[snake_writer_iterator], SNAKE};
							if(snake_writer_iterator == snake_size+16'd1)
							begin
								rect_write_nxt = {snake_register[snake_writer_iterator], NULL};
								snake_register_nxt[snake_writer_iterator] = 0;
							end

							if(snake_writer_iterator == SNAKE_REG_SIZE) snake_writer_iterator_nxt = 0;
							else snake_writer_iterator_nxt = snake_writer_iterator + 16'd1;
						end

					COLLISION_READ:
						begin
							state_nxt = COLLISION_CHECK;
							rect_read_out_nxt = snake_register[0];
						end

					COLLISION_CHECK:
						begin
							case(rect_read_in)
								SNAKE:
									state_nxt = GAME_OVER;
								SNACK:
									state_nxt = SNAKE_GROW;
								ROCK:
									state_nxt = GAME_OVER;
								default:
									state_nxt = SNAKE_DRAWING;
							endcase
						end

					SNAKE_GROW:
						begin
							snake_size_nxt = snake_size + 5'd1;
							state_nxt = SNACK_GENERATE;
							snake_writer_iterator_nxt = 0;
							score_nxt = score_out + (difficulty_level*16'd10)/2;
							if (snake_speed <= 20000000/difficulty_level) snake_speed_nxt = snake_speed;
							else 	snake_speed_nxt = snake_speed - difficulty_level*1000000;
						end

					GAME_OVER:
						begin
							if(rst) state_nxt = INIT;
							else if(game_restart == 1) state_nxt = INIT;
							else state_nxt = GAME_OVER;
							game_over_nxt = 1;
						end

					SNACK_GENERATE:
						begin
							state_nxt = SNACK_CHECK_READ;
							for(i = 0; i <= 31; i=i+1)
								{snack_gen_reg_x_nxt,snack_gen_reg_y_nxt} ={snack_gen_reg_x_nxt+snake_register[i][4:0],snack_gen_reg_y_nxt+snake_register[i][20:16]} ;
						end

					SNACK_CHECK_READ:
						begin
							state_nxt = SNACK_CHECK_WRITE;
							rect_read_out_nxt = {11'b0, snack_gen_reg_x, 11'b0, snack_gen_reg_y};
							//		rect_read_out_nxt[20:16] = snack_gen_reg_x;
							//		rect_read_out_nxt[4:0] = snack_gen_reg_y;
						end

					SNACK_CHECK_WRITE:
						begin
							state_nxt = SNACK_CHECK_READ;
							if(rect_read_in != NULL)
								begin
									{snack_gen_reg_x_nxt,snack_gen_reg_y_nxt} =  {snack_gen_reg_x+snake_register[2][4:0],snack_gen_reg_y+snake_register[2][20:16]};
								end
							else
								begin
									rect_write_nxt = 32'b0;
									rect_write_nxt[24:20] = snack_gen_reg_x;
									rect_write_nxt[8:4] = snack_gen_reg_y;
									rect_write_nxt[3:0] = SNACK;
									state_nxt = SNAKE_DRAWING;
								end
							//TODO snack on snake checking
						end
					MENU_INTERRUPT:
						begin
							if(menu_interrupt == 0)state_nxt = SNAKE_DRAWING;
							else state_nxt = MENU_INTERRUPT;
							snake_moving_iterator_nxt = snake_moving_iterator;
						end			
				endcase

			if(rst) state_nxt = WAIT_FOR_START;	
		end
   			
   always@(posedge clk)
      begin
				snake_writer_iterator <= snake_writer_iterator_nxt;
				snake_moving_iterator <= snake_moving_iterator_nxt;
				snake_size <= snake_size_nxt;
				state <= state_nxt;
				rect_write <= rect_write_nxt;
				rect_read_out <= rect_read_out_nxt;
				snack_gen_reg_y <= snack_gen_reg_y_nxt; 
				snack_gen_reg_x<= snack_gen_reg_x_nxt; 
				snake_speed <= snake_speed_nxt;
				score_out <= score_nxt;
				game_over <= game_over_nxt;
      end
        
genvar X;		
	generate
			begin
			for (X = 0; X <= SNAKE_REG_SIZE; X = X+1)		
				begin
					always@(posedge clk)
						begin
							snake_register[X] <= snake_register_nxt[X];
						end	
				end
			end	
	endgenerate	 
	
	
	/*
     //DEBUG DISPLAY
	reg [3:0] hex3, hex2, hex1, hex0;  // hex digits
    wire [3:0] dp_in;             // 4 decimal points
	wire [31:0] rx;
	
	assign rx = snake_register[debug_keys];
	always@(*)
	begin
		if(debug_keys == 5'b11111) //State debug
			begin
				hex3 = 0;
				hex2 = 0;
				hex1 = 0;
				hex0 = state;
			end
		else if(debug_keys == 5'b11110)	//GRID REGISTER READ DEBUG
			begin
				hex3 = 0;
				hex2 = 0;
				hex1 = 0;
				hex0 = rect_read_in;
			end
		else if(debug_keys == 5'b11100)	
			begin
				{hex3, hex2, hex1, hex0} = {3'b0, snack_gen_reg_x, 3'b0, snack_gen_reg_y}; //SNACK GENERATION DEBUG
			end			
		else if(debug_keys == 5'b11101)	
			begin
				{hex3, hex2, hex1, hex0} = snake_speed/1000000; //SNAKE SPEED
			end
		else if(debug_keys == 5'b11001)	
			begin
				{hex3, hex2, hex1, hex0} = {snake_size}; //SNAKE_SIZE
			end
		else if(debug_keys == 5'b10101)	
			begin
				{hex3, hex2, hex1, hex0} = {r_data}; //r_read 
			end
		else if(debug_keys == 5'b00101)	
			begin
				{hex3, hex2, hex1, hex0} = iterator_debug; //r_read 
			end									
		else		
	// 	{hex3, hex2, hex1, hex0} = {rx[23:16],rx[7:0]};
			{hex3, hex2, hex1, hex0} = 16'hFFFF;
	end

   // constant declaration
   // refreshing rate around 800 Hz (50 MHz/2^16)
   localparam N = 18;
   // internal signal declaration
   reg [N-1:0] q_reg;
   wire [N-1:0] q_next;
   reg [3:0] hex_in;
   reg dp;

   // N-bit counter
   // register
   always @(posedge clk, posedge rst)
      if (rst)
         q_reg <= 0;
      else
         q_reg <= q_next;

   // next-state logic
   assign q_next = q_reg + 1;

   // 2 MSBs of counter to control 4-to-1 multiplexing
   // and to generate active-low enable signal
   always @*
      case (q_reg[N-1:N-2])
         2'b00:
            begin
               an =  4'b1110;
               hex_in = hex0;
               dp = dp_in[0];
            end
         2'b01:
            begin
               an =  4'b1101;
               hex_in = hex1;
               dp = dp_in[1];
            end
         2'b10:
            begin
               an =  4'b1011;
               hex_in = hex2;
               dp = dp_in[2];
            end
         default:
            begin
               an =  4'b0111;
               hex_in = hex3;
               dp = dp_in[3];
            end
       endcase

   // hex to seven-segment led display
   always @*
   begin
      case(hex_in)
         4'h0: sseg[6:0] = 7'b0000001;
         4'h1: sseg[6:0] = 7'b1001111;
         4'h2: sseg[6:0] = 7'b0010010;
         4'h3: sseg[6:0] = 7'b0000110;
         4'h4: sseg[6:0] = 7'b1001100;
         4'h5: sseg[6:0] = 7'b0100100;
         4'h6: sseg[6:0] = 7'b0100000;
         4'h7: sseg[6:0] = 7'b0001111;
         4'h8: sseg[6:0] = 7'b0000000;
         4'h9: sseg[6:0] = 7'b0000100;
         4'ha: sseg[6:0] = 7'b0001000;
         4'hb: sseg[6:0] = 7'b1100000;
         4'hc: sseg[6:0] = 7'b0110001;
         4'hd: sseg[6:0] = 7'b1000010;
         4'he: sseg[6:0] = 7'b0110000;
         default: sseg[6:0] = 7'b0111000;  //4'hf
     endcase
   end


	 
    
    
   */
endmodule
